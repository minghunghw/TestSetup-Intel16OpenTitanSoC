#############################################################################################
## Intel Confidential                                                                      ##
#############################################################################################
## Copyright 2022 Intel Corporation. The information contained herein is the proprietary   ##
## and confidential information of Intel or its licensors, and is supplied subject to, and ##
## may be used only in accordance with, previously executed agreements with Intel.         ##
## EXCEPT AS MAY OTHERWISE BE AGREED IN WRITING: (1) ALL MATERIALS FURNISHED BY INTEL      ##
## HEREUNDER ARE PROVIDED "AS IS" WITHOUT WARRANTY OF ANY KIND; (2) INTEL SPECIFICALLY     ##
## DISCLAIMS ANY WARRANTY OF NONINFRINGEMENT, FITNESS FOR A PARTICULAR PURPOSE OR          ##
## MERCHANTABILITY; AND (3) INTEL WILL NOT BE LIABLE FOR ANY COSTS OF PROCUREMENT OF       ##
## SUBSTITUTES, LOSS OF PROFITS, INTERRUPTION OF BUSINESS, OR FOR ANY OTHER SPECIAL,       ##
## CONSEQUENTIAL OR INCIDENTAL DAMAGES, HOWEVER CAUSED, WHETHER FOR BREACH OF WARRANTY,    ##
## CONTRACT, TORT, NEGLIGENCE, STRICT LIABILITY OR OTHERWISE.                              ##
#############################################################################################
#############################################################################################
##                                                                                         ##
##  Vendor:                Intel Corporation                                               ##
##  Product:               ip224uhdlp1p11rf                                                ##
##  Version:               r1.0.1                                                          ##
##  Technology:            p1222.4                                                         ##
##  Celltype:              MemoryIP                                                        ##
##  IP Owner:              Intel CMO                                                       ##
##  Creation Time:         Wed Sep 14 2022 15:14:42                                        ##
##  Memory Name:           ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p0d0a1m1h                  ##
##  Memory Name Generated: ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p0d0a1m1h                  ##
##                                                                                         ##
#############################################################################################

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
SITE ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p0d0a1m1h
  SIZE 134.396 by 65.7 ;
  SYMMETRY X Y ;
  CLASS CORE ;
END ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p0d0a1m1h


MACRO ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p0d0a1m1h
     FOREIGN ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p0d0a1m1h 0.00 0.00 ;
     ORIGIN 0.00 0.00 ;
     SIZE 134.396 by 65.7 ;
     SYMMETRY X Y ;
     CLASS BLOCK ;
     SITE ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p0d0a1m1h ;
     PIN adr[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 73.7555 37.004 74.9455 37.08 ;
          END
     END adr[0]
     PIN adr[10]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 61.5735 37.3 62.525 37.376 ;
          END
     END adr[10]
     PIN adr[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 73.3605 35.884 74.3475 35.96 ;
          END
     END adr[1]
     PIN adr[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 73.186 34.928 74.36 35.004 ;
          END
     END adr[2]
     PIN adr[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 74.44 34.928 75.39 35.004 ;
          END
     END adr[3]
     PIN adr[4]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 58.641 27.04 59.598 27.116 ;
          END
     END adr[4]
     PIN adr[5]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 59.9225 32.406 60.862 32.462 ;
          END
     END adr[5]
     PIN adr[6]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 59.362 28.306 60.4255 28.382 ;
          END
     END adr[6]
     PIN adr[7]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 58.988 28.456 60.337 28.532 ;
          END
     END adr[7]
     PIN adr[8]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 61.291 35.884 62.2155 35.96 ;
          END
     END adr[8]
     PIN adr[9]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 61.303 37.004 62.433 37.08 ;
          END
     END adr[9]
     PIN clkbyp
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 70.363 32.406 71.2155 32.462 ;
          END
     END clkbyp
     PIN din[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 64.268 65.283 64.376 ;
          END
     END din[0]
     PIN din[10]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 48.068 65.283 48.176 ;
          END
     END din[10]
     PIN din[11]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 46.448 65.283 46.556 ;
          END
     END din[11]
     PIN din[12]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 44.828 65.283 44.936 ;
          END
     END din[12]
     PIN din[13]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 43.208 65.283 43.316 ;
          END
     END din[13]
     PIN din[14]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 41.588 65.283 41.696 ;
          END
     END din[14]
     PIN din[15]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 39.968 65.283 40.076 ;
          END
     END din[15]
     PIN din[16]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 25.748 65.283 25.856 ;
          END
     END din[16]
     PIN din[17]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 24.128 65.283 24.236 ;
          END
     END din[17]
     PIN din[18]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 22.508 65.283 22.616 ;
          END
     END din[18]
     PIN din[19]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 20.888 65.283 20.996 ;
          END
     END din[19]
     PIN din[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 62.648 65.283 62.756 ;
          END
     END din[1]
     PIN din[20]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 19.268 65.283 19.376 ;
          END
     END din[20]
     PIN din[21]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 17.648 65.283 17.756 ;
          END
     END din[21]
     PIN din[22]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 16.028 65.283 16.136 ;
          END
     END din[22]
     PIN din[23]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 14.408 65.283 14.516 ;
          END
     END din[23]
     PIN din[24]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 12.788 65.283 12.896 ;
          END
     END din[24]
     PIN din[25]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 11.168 65.283 11.276 ;
          END
     END din[25]
     PIN din[26]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 9.548 65.283 9.656 ;
          END
     END din[26]
     PIN din[27]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 7.928 65.283 8.036 ;
          END
     END din[27]
     PIN din[28]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 6.308 65.283 6.416 ;
          END
     END din[28]
     PIN din[29]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 4.688 65.283 4.796 ;
          END
     END din[29]
     PIN din[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 61.028 65.283 61.136 ;
          END
     END din[2]
     PIN din[30]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 3.068 65.283 3.176 ;
          END
     END din[30]
     PIN din[31]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 1.448 65.283 1.556 ;
          END
     END din[31]
     PIN din[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 59.408 65.283 59.516 ;
          END
     END din[3]
     PIN din[4]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 57.788 65.283 57.896 ;
          END
     END din[4]
     PIN din[5]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 56.168 65.283 56.276 ;
          END
     END din[5]
     PIN din[6]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 54.548 65.283 54.656 ;
          END
     END din[6]
     PIN din[7]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 52.928 65.283 53.036 ;
          END
     END din[7]
     PIN din[8]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 51.308 65.283 51.416 ;
          END
     END din[8]
     PIN din[9]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.9205 49.688 65.283 49.796 ;
          END
     END din[9]
     PIN fwen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 74.0155 31.57 75.702 31.626 ;
          END
     END fwen
     PIN mc[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 60.84 34.204 61.879 34.28 ;
          END
     END mc[0]
     PIN mc[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 58.62 35.62 59.848 35.696 ;
          END
     END mc[1]
     PIN mc[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 59.979 35.62 61.121 35.696 ;
          END
     END mc[2]
     PIN mcen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 60.0765 35.884 61.013 35.96 ;
          END
     END mcen
     PIN q[0]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 64.268 67.7695 64.376 ;
          END
     END q[0]
     PIN q[10]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 48.068 67.7695 48.176 ;
          END
     END q[10]
     PIN q[11]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 46.448 67.7695 46.556 ;
          END
     END q[11]
     PIN q[12]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 44.828 67.7695 44.936 ;
          END
     END q[12]
     PIN q[13]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 43.208 67.7695 43.316 ;
          END
     END q[13]
     PIN q[14]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 41.588 67.7695 41.696 ;
          END
     END q[14]
     PIN q[15]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 39.968 67.7695 40.076 ;
          END
     END q[15]
     PIN q[16]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 25.748 67.7695 25.856 ;
          END
     END q[16]
     PIN q[17]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 24.128 67.7695 24.236 ;
          END
     END q[17]
     PIN q[18]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 22.508 67.7695 22.616 ;
          END
     END q[18]
     PIN q[19]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 20.888 67.7695 20.996 ;
          END
     END q[19]
     PIN q[1]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 62.648 67.7695 62.756 ;
          END
     END q[1]
     PIN q[20]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 19.268 67.7695 19.376 ;
          END
     END q[20]
     PIN q[21]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 17.648 67.7695 17.756 ;
          END
     END q[21]
     PIN q[22]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 16.028 67.7695 16.136 ;
          END
     END q[22]
     PIN q[23]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 14.408 67.7695 14.516 ;
          END
     END q[23]
     PIN q[24]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 12.788 67.7695 12.896 ;
          END
     END q[24]
     PIN q[25]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 11.168 67.7695 11.276 ;
          END
     END q[25]
     PIN q[26]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 9.548 67.7695 9.656 ;
          END
     END q[26]
     PIN q[27]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 7.928 67.7695 8.036 ;
          END
     END q[27]
     PIN q[28]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 6.308 67.7695 6.416 ;
          END
     END q[28]
     PIN q[29]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 4.688 67.7695 4.796 ;
          END
     END q[29]
     PIN q[2]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 61.028 67.7695 61.136 ;
          END
     END q[2]
     PIN q[30]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 3.068 67.7695 3.176 ;
          END
     END q[30]
     PIN q[31]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 1.448 67.7695 1.556 ;
          END
     END q[31]
     PIN q[3]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 59.408 67.7695 59.516 ;
          END
     END q[3]
     PIN q[4]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 57.788 67.7695 57.896 ;
          END
     END q[4]
     PIN q[5]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 56.168 67.7695 56.276 ;
          END
     END q[5]
     PIN q[6]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 54.548 67.7695 54.656 ;
          END
     END q[6]
     PIN q[7]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 52.928 67.7695 53.036 ;
          END
     END q[7]
     PIN q[8]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 51.308 67.7695 51.416 ;
          END
     END q[8]
     PIN q[9]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 65.8185 49.688 67.7695 49.796 ;
          END
     END q[9]
     PIN ren
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 69.746 31.57 70.6515 31.626 ;
          END
     END ren
     PIN wa[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 72.308 33.938 73.2725 33.994 ;
          END
     END wa[0]
     PIN wa[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 71.0955 33.938 72.126 33.994 ;
          END
     END wa[1]
     PIN wen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 71.21 31.57 72.098 31.626 ;
          END
     END wen
     PIN wpulse[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 73.835 30.004 74.8205 30.08 ;
          END
     END wpulse[0]
     PIN wpulse[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 69.3545 29.28 70.398 29.356 ;
          END
     END wpulse[1]
     PIN wpulseen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 70.1605 30.004 71.047 30.08 ;
          END
     END wpulseen
     PIN clk
     DIRECTION input ;
          USE CLOCK ;
          PORT
               LAYER m4 ;
               RECT 67.8205 32.406 68.8525 32.462 ;
          END
     END clk
     PIN vddp
     SHAPE ABUTMENT ;
     DIRECTION input ;
          USE POWER ;
          PORT
               LAYER m4 ;
               RECT 0.48 0.958 61.218 1.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 1.846 57.036 1.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 10.678 61.218 10.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 11.566 57.036 11.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 12.298 61.218 12.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.186 57.036 13.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.918 61.218 13.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 14.806 57.036 14.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 15.538 61.218 15.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 16.426 57.036 16.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 17.158 61.218 17.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.046 57.036 18.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.778 61.218 18.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 19.666 57.036 19.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 2.578 61.218 2.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 20.398 61.218 20.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 21.286 57.036 21.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 22.018 61.218 22.094 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 22.906 57.036 22.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 23.638 61.218 23.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 24.526 57.036 24.602 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 25.258 61.218 25.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 26.146 57.036 26.222 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 3.466 57.036 3.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 39.478 61.218 39.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 4.198 61.218 4.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 40.366 57.036 40.442 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 41.098 61.218 41.174 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 41.986 57.036 42.062 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 42.718 61.218 42.794 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 43.606 57.036 43.682 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 44.338 61.218 44.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 45.226 57.036 45.302 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 45.958 61.218 46.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 46.846 57.036 46.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 47.578 61.218 47.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 48.466 57.036 48.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 49.198 61.218 49.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.086 57.036 5.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.818 61.218 5.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 50.086 57.036 50.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 50.818 61.218 50.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 51.706 57.036 51.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 52.438 61.218 52.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 53.326 57.036 53.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 54.058 61.218 54.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 54.946 57.036 55.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 55.678 61.218 55.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 56.566 57.036 56.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 57.298 61.218 57.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 58.186 57.036 58.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 58.918 61.218 58.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 59.806 57.036 59.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 6.706 57.036 6.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 60.538 61.218 60.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 61.426 57.036 61.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 62.158 61.218 62.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 63.046 57.036 63.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 63.778 61.218 63.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 64.666 57.036 64.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 7.438 61.218 7.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 8.326 57.036 8.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 9.058 61.218 9.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 9.946 57.036 10.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 28.028 57.208 28.104 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 28.588 133.78 28.664 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 28.984 133.78 29.06 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 29.28 57.208 29.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 30.004 57.208 30.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 31.072 56.56 31.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 31.57 57.208 31.626 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 32.406 57.208 32.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 33.324 56.56 33.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 34.336 133.78 34.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 35.06 133.78 35.136 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 35.356 133.78 35.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 35.752 133.78 35.828 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 36.312 133.78 36.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 38.256 133.78 38.364 ;
          END
          PORT
               LAYER m4 ;
               RECT 1.264 29.712 56.56 29.82 ;
          END
          PORT
               LAYER m4 ;
               RECT 1.264 30.268 56.56 30.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 1.264 34.04 56.56 34.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 1.264 34.596 56.56 34.704 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 26.644 77.148 26.72 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 27.896 77.148 27.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 29.412 77.148 29.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 38.98 77.148 39.056 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.317 30.004 70.0805 30.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.348 34.05 77.1075 34.126 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 1.324 77.033 1.4 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 11.044 77.033 11.12 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 12.664 77.033 12.74 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 14.284 77.033 14.36 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 15.904 77.033 15.98 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 17.524 77.033 17.6 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 19.144 77.033 19.22 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 2.944 77.033 3.02 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 20.764 77.033 20.84 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 22.384 77.033 22.46 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 24.004 77.033 24.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 25.624 77.033 25.7 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 39.844 77.033 39.92 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 4.564 77.033 4.64 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 41.464 77.033 41.54 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 43.084 77.033 43.16 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 44.704 77.033 44.78 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 46.324 77.033 46.4 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 47.944 77.033 48.02 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 49.564 77.033 49.64 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 51.184 77.033 51.26 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 52.804 77.033 52.88 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 54.424 77.033 54.5 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 56.044 77.033 56.12 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 57.664 77.033 57.74 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 59.284 77.033 59.36 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 6.184 77.033 6.26 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 60.904 77.033 60.98 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 62.524 77.033 62.6 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 64.144 77.033 64.22 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 7.804 77.033 7.88 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.503 9.424 77.033 9.5 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 1.08 73.295 1.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 10.8 73.295 10.876 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 12.42 73.295 12.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 14.04 73.295 14.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 15.66 73.295 15.736 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 17.28 73.295 17.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 18.9 73.295 18.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 2.7 73.295 2.776 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 20.52 73.295 20.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 22.14 73.295 22.216 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 23.76 73.295 23.836 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 25.38 73.295 25.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 39.6 73.295 39.676 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 4.32 73.295 4.396 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 41.22 73.295 41.296 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 42.84 73.295 42.916 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 44.46 73.295 44.536 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 46.08 73.295 46.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 47.7 73.295 47.776 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 49.32 73.295 49.396 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 5.94 73.295 6.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 50.94 73.295 51.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 52.56 73.295 52.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 54.18 73.295 54.256 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 55.8 73.295 55.876 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 57.42 73.295 57.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 59.04 73.295 59.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 60.66 73.295 60.736 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 62.28 73.295 62.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 63.9 73.295 63.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 7.56 73.295 7.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 61.142 9.18 73.295 9.256 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 0.958 133.916 1.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 10.678 133.916 10.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 12.298 133.916 12.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 13.918 133.916 13.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 15.538 133.916 15.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 17.158 133.916 17.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 18.778 133.916 18.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 2.578 133.916 2.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 20.398 133.916 20.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 22.018 133.916 22.094 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 23.638 133.916 23.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 25.258 133.916 25.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 39.478 133.916 39.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 4.198 133.916 4.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 41.098 133.916 41.174 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 42.718 133.916 42.794 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 44.338 133.916 44.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 45.958 133.916 46.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 47.578 133.916 47.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 49.198 133.916 49.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 5.818 133.916 5.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 50.818 133.916 50.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 52.438 133.916 52.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 54.058 133.916 54.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 55.678 133.916 55.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 57.298 133.916 57.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 58.918 133.916 58.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 60.538 133.916 60.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 62.158 133.916 62.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 63.778 133.916 63.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 7.438 133.916 7.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.219 9.058 133.916 9.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 28.028 133.78 28.104 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 30.004 133.78 30.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 31.57 133.78 31.626 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 32.406 133.78 32.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.228 29.28 133.78 29.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 1.846 133.916 1.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 11.566 133.916 11.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 13.186 133.916 13.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 14.806 133.916 14.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 16.426 133.916 16.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 18.046 133.916 18.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 19.666 133.916 19.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 21.286 133.916 21.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 22.906 133.916 22.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 24.526 133.916 24.602 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 26.146 133.916 26.222 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 3.466 133.916 3.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 40.366 133.916 40.442 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 41.986 133.916 42.062 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 43.606 133.916 43.682 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 45.226 133.916 45.302 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 46.846 133.916 46.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 48.466 133.916 48.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 5.086 133.916 5.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 50.086 133.916 50.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 51.706 133.916 51.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 53.326 133.916 53.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 54.946 133.916 55.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 56.566 133.916 56.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 58.186 133.916 58.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 59.806 133.916 59.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 6.706 133.916 6.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 61.426 133.916 61.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 63.046 133.916 63.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 64.666 133.916 64.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 8.326 133.916 8.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.293 9.946 133.916 10.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.836 29.712 133.132 29.82 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.836 30.268 133.132 30.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.836 31.072 133.78 31.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.836 33.324 133.78 33.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.836 34.04 133.132 34.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.836 34.596 133.78 34.704 ;
          END
     END vddp
     PIN vss
     SHAPE ABUTMENT ;
     DIRECTION inout ;
          USE GROUND ;
          PORT
               LAYER m4 ;
               RECT 0.48 0.592 77.1815 0.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 10.312 77.1815 10.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 11.932 77.1815 12.008 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.552 77.1815 13.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 15.172 77.1815 15.248 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 16.792 77.1815 16.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.412 77.1815 18.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 2.212 77.1815 2.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 20.032 77.1815 20.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 21.652 77.1815 21.728 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 23.272 77.1815 23.348 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 24.892 77.1815 24.968 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 26.512 133.916 26.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 3.832 77.1815 3.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 39.112 133.916 39.188 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 40.732 77.1815 40.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 42.352 77.1815 42.428 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 43.972 77.1815 44.048 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 45.592 77.1815 45.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 47.212 77.1815 47.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 48.832 77.1815 48.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.452 77.1815 5.528 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 50.452 77.1815 50.528 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 52.072 77.1815 52.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 53.692 77.1815 53.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 55.312 77.1815 55.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 56.932 77.1815 57.008 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 58.552 77.1815 58.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 60.172 77.1815 60.248 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 61.792 77.1815 61.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 63.412 77.1815 63.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 65.032 77.1815 65.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 7.072 77.1815 7.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 8.692 77.1815 8.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 27.172 77.836 27.28 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 27.468 77.836 27.576 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 29.544 77.836 29.652 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 30.566 57.208 30.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 30.982 77.836 31.026 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 32.08 77.836 32.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 33.414 77.836 33.458 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 33.83 57.208 33.874 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 34.764 77.836 34.872 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 36.84 77.836 36.948 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 37.136 77.836 37.244 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 37.96 77.836 38.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 38.552 77.836 38.66 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.208 30.554 77.0235 30.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.35 33.836 77.1075 33.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 1.602 76.9585 1.678 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 11.322 76.9585 11.398 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 12.942 76.9585 13.018 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 14.562 76.9585 14.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 16.182 76.9585 16.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 17.802 76.9585 17.878 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 19.422 76.9585 19.498 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 21.042 76.9585 21.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 22.662 76.9585 22.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 24.282 76.9585 24.358 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 25.902 76.9585 25.978 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 3.222 76.9585 3.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 4.842 76.9585 4.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 40.122 76.9585 40.198 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 41.742 76.9585 41.818 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 43.362 76.9585 43.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 44.982 76.9585 45.058 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 46.602 76.9585 46.678 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 48.222 76.9585 48.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 49.842 76.9585 49.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 51.462 76.9585 51.538 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 53.082 76.9585 53.158 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 54.702 76.9585 54.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 56.322 76.9585 56.398 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 57.942 76.9585 58.018 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 59.562 76.9585 59.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 6.462 76.9585 6.538 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 61.182 76.9585 61.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 62.802 76.9585 62.878 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 64.422 76.9585 64.498 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 8.082 76.9585 8.158 ;
          END
          PORT
               LAYER m4 ;
               RECT 59.9355 9.702 76.9585 9.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 0.592 133.916 0.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 10.312 133.916 10.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 11.932 133.916 12.008 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 13.552 133.916 13.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 15.172 133.916 15.248 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 16.792 133.916 16.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 18.412 133.916 18.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 2.212 133.916 2.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 20.032 133.916 20.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 21.652 133.916 21.728 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 23.272 133.916 23.348 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 24.892 133.916 24.968 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 3.832 133.916 3.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 40.732 133.916 40.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 42.352 133.916 42.428 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 43.972 133.916 44.048 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 45.592 133.916 45.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 47.212 133.916 47.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 48.832 133.916 48.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 5.452 133.916 5.528 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 50.452 133.916 50.528 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 52.072 133.916 52.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 53.692 133.916 53.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 55.312 133.916 55.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 56.932 133.916 57.008 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 58.552 133.916 58.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 60.172 133.916 60.248 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 61.792 133.916 61.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 63.412 133.916 63.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 65.032 133.916 65.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 7.072 133.916 7.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.188 8.692 133.916 8.768 ;
          END
     END vss
     OBS
          LAYER m1 SPACING 0 ;
               RECT 0.248 0.198 134.148 65.502 ;
          LAYER m2 SPACING 0 ;
               RECT 0.32 0.268 134.076 65.432 ;
          LAYER m3 SPACING 0 ;
               RECT 0.342 0.24 134.054 65.46 ;
          LAYER m4 SPACING 0 ;
               RECT 0.32 0.31 134.076 65.34 ;
     END
END ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p0d0a1m1h
END LIBRARY
