#############################################################################################
## Intel Confidential                                                                      ##
#############################################################################################
## Copyright 2022 Intel Corporation. The information contained herein is the proprietary   ##
## and confidential information of Intel or its licensors, and is supplied subject to, and ##
## may be used only in accordance with, previously executed agreements with Intel.         ##
## EXCEPT AS MAY OTHERWISE BE AGREED IN WRITING: (1) ALL MATERIALS FURNISHED BY INTEL      ##
## HEREUNDER ARE PROVIDED "AS IS" WITHOUT WARRANTY OF ANY KIND; (2) INTEL SPECIFICALLY     ##
## DISCLAIMS ANY WARRANTY OF NONINFRINGEMENT, FITNESS FOR A PARTICULAR PURPOSE OR          ##
## MERCHANTABILITY; AND (3) INTEL WILL NOT BE LIABLE FOR ANY COSTS OF PROCUREMENT OF       ##
## SUBSTITUTES, LOSS OF PROFITS, INTERRUPTION OF BUSINESS, OR FOR ANY OTHER SPECIAL,       ##
## CONSEQUENTIAL OR INCIDENTAL DAMAGES, HOWEVER CAUSED, WHETHER FOR BREACH OF WARRANTY,    ##
## CONTRACT, TORT, NEGLIGENCE, STRICT LIABILITY OR OTHERWISE.                              ##
#############################################################################################
#############################################################################################
##                                                                                         ##
##  Vendor:                Intel Corporation                                               ##
##  Product:               ip224uhdlp1p11rf                                                ##
##  Version:               r1.0.1                                                          ##
##  Technology:            p1222.4                                                         ##
##  Celltype:              MemoryIP                                                        ##
##  IP Owner:              Intel CMO                                                       ##
##  Creation Time:         Wed Sep 14 2022 15:16:23                                        ##
##  Memory Name:           ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p1d0a1m1h                  ##
##  Memory Name Generated: ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p1d0a1m1h                  ##
##                                                                                         ##
#############################################################################################

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
SITE ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p1d0a1m1h
  SIZE 138.5 by 65.7 ;
  SYMMETRY X Y ;
  CLASS CORE ;
END ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p1d0a1m1h


MACRO ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p1d0a1m1h
     FOREIGN ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p1d0a1m1h 0.00 0.00 ;
     ORIGIN 0.00 0.00 ;
     SIZE 138.5 by 65.7 ;
     SYMMETRY X Y ;
     CLASS BLOCK ;
     SITE ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p1d0a1m1h ;
     PIN adr[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 75.8075 37.004 76.9975 37.08 ;
          END
     END adr[0]
     PIN adr[10]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.6255 37.3 64.577 37.376 ;
          END
     END adr[10]
     PIN adr[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 75.4125 35.884 76.3995 35.96 ;
          END
     END adr[1]
     PIN adr[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 75.238 34.928 76.412 35.004 ;
          END
     END adr[2]
     PIN adr[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 76.492 34.928 77.654 35.004 ;
          END
     END adr[3]
     PIN adr[4]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 60.693 27.04 61.65 27.116 ;
          END
     END adr[4]
     PIN adr[5]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 61.9745 32.406 62.914 32.462 ;
          END
     END adr[5]
     PIN adr[6]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 60.656 28.306 62.037 28.382 ;
          END
     END adr[6]
     PIN adr[7]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 61.0805 28.456 62.389 28.532 ;
          END
     END adr[7]
     PIN adr[8]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.343 35.884 64.2675 35.96 ;
          END
     END adr[8]
     PIN adr[9]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 63.355 37.004 64.485 37.08 ;
          END
     END adr[9]
     PIN bc1
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 75.4925 35.62 76.5565 35.696 ;
          END
     END bc1
     PIN bc2
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 76.412 33.938 77.5515 33.994 ;
          END
     END bc2
     PIN clkbyp
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 72.415 32.406 73.2675 32.462 ;
          END
     END clkbyp
     PIN deepslp
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 76.916 32.406 77.91 32.462 ;
          END
     END deepslp
     PIN din[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 64.268 67.1525 64.376 ;
          END
     END din[0]
     PIN din[10]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 48.068 67.1525 48.176 ;
          END
     END din[10]
     PIN din[11]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 46.448 67.1525 46.556 ;
          END
     END din[11]
     PIN din[12]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 44.828 67.1525 44.936 ;
          END
     END din[12]
     PIN din[13]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 43.208 67.1525 43.316 ;
          END
     END din[13]
     PIN din[14]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 41.588 67.1525 41.696 ;
          END
     END din[14]
     PIN din[15]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 39.968 67.1525 40.076 ;
          END
     END din[15]
     PIN din[16]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 25.748 67.1525 25.856 ;
          END
     END din[16]
     PIN din[17]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 24.128 67.1525 24.236 ;
          END
     END din[17]
     PIN din[18]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 22.508 67.1525 22.616 ;
          END
     END din[18]
     PIN din[19]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 20.888 67.1525 20.996 ;
          END
     END din[19]
     PIN din[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 62.648 67.1525 62.756 ;
          END
     END din[1]
     PIN din[20]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 19.268 67.1525 19.376 ;
          END
     END din[20]
     PIN din[21]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 17.648 67.1525 17.756 ;
          END
     END din[21]
     PIN din[22]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 16.028 67.1525 16.136 ;
          END
     END din[22]
     PIN din[23]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 14.408 67.1525 14.516 ;
          END
     END din[23]
     PIN din[24]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 12.788 67.1525 12.896 ;
          END
     END din[24]
     PIN din[25]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 11.168 67.1525 11.276 ;
          END
     END din[25]
     PIN din[26]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 9.548 67.1525 9.656 ;
          END
     END din[26]
     PIN din[27]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 7.928 67.1525 8.036 ;
          END
     END din[27]
     PIN din[28]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 6.308 67.1525 6.416 ;
          END
     END din[28]
     PIN din[29]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 4.688 67.1525 4.796 ;
          END
     END din[29]
     PIN din[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 61.028 67.1525 61.136 ;
          END
     END din[2]
     PIN din[30]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 3.068 67.1525 3.176 ;
          END
     END din[30]
     PIN din[31]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 1.448 67.1525 1.556 ;
          END
     END din[31]
     PIN din[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 59.408 67.1525 59.516 ;
          END
     END din[3]
     PIN din[4]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 57.788 67.1525 57.896 ;
          END
     END din[4]
     PIN din[5]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 56.168 67.1525 56.276 ;
          END
     END din[5]
     PIN din[6]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 54.548 67.1525 54.656 ;
          END
     END din[6]
     PIN din[7]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 52.928 67.1525 53.036 ;
          END
     END din[7]
     PIN din[8]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 51.308 67.1525 51.416 ;
          END
     END din[8]
     PIN din[9]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 64.658 49.688 67.1525 49.796 ;
          END
     END din[9]
     PIN fwen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 76.0675 31.57 77.022 31.626 ;
          END
     END fwen
     PIN mc[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 62.892 34.204 63.931 34.28 ;
          END
     END mc[0]
     PIN mc[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 60.672 35.62 61.9 35.696 ;
          END
     END mc[1]
     PIN mc[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 62.031 35.62 63.173 35.696 ;
          END
     END mc[2]
     PIN mcen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 62.1285 35.884 63.065 35.96 ;
          END
     END mcen
     PIN mpr
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 74.773 31.57 75.709 31.626 ;
          END
     END mpr
     PIN q[0]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 64.268 69.3865 64.376 ;
          END
     END q[0]
     PIN q[10]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 48.068 69.3865 48.176 ;
          END
     END q[10]
     PIN q[11]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 46.448 69.3865 46.556 ;
          END
     END q[11]
     PIN q[12]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 44.828 69.3865 44.936 ;
          END
     END q[12]
     PIN q[13]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 43.208 69.3865 43.316 ;
          END
     END q[13]
     PIN q[14]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 41.588 69.3865 41.696 ;
          END
     END q[14]
     PIN q[15]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 39.968 69.3865 40.076 ;
          END
     END q[15]
     PIN q[16]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 25.748 69.3865 25.856 ;
          END
     END q[16]
     PIN q[17]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 24.128 69.3865 24.236 ;
          END
     END q[17]
     PIN q[18]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 22.508 69.3865 22.616 ;
          END
     END q[18]
     PIN q[19]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 20.888 69.3865 20.996 ;
          END
     END q[19]
     PIN q[1]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 62.648 69.3865 62.756 ;
          END
     END q[1]
     PIN q[20]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 19.268 69.3865 19.376 ;
          END
     END q[20]
     PIN q[21]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 17.648 69.3865 17.756 ;
          END
     END q[21]
     PIN q[22]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 16.028 69.3865 16.136 ;
          END
     END q[22]
     PIN q[23]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 14.408 69.3865 14.516 ;
          END
     END q[23]
     PIN q[24]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 12.788 69.3865 12.896 ;
          END
     END q[24]
     PIN q[25]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 11.168 69.3865 11.276 ;
          END
     END q[25]
     PIN q[26]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 9.548 69.3865 9.656 ;
          END
     END q[26]
     PIN q[27]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 7.928 69.3865 8.036 ;
          END
     END q[27]
     PIN q[28]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 6.308 69.3865 6.416 ;
          END
     END q[28]
     PIN q[29]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 4.688 69.3865 4.796 ;
          END
     END q[29]
     PIN q[2]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 61.028 69.3865 61.136 ;
          END
     END q[2]
     PIN q[30]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 3.068 69.3865 3.176 ;
          END
     END q[30]
     PIN q[31]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 1.448 69.3865 1.556 ;
          END
     END q[31]
     PIN q[3]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 59.408 69.3865 59.516 ;
          END
     END q[3]
     PIN q[4]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 57.788 69.3865 57.896 ;
          END
     END q[4]
     PIN q[5]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 56.168 69.3865 56.276 ;
          END
     END q[5]
     PIN q[6]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 54.548 69.3865 54.656 ;
          END
     END q[6]
     PIN q[7]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 52.928 69.3865 53.036 ;
          END
     END q[7]
     PIN q[8]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 51.308 69.3865 51.416 ;
          END
     END q[8]
     PIN q[9]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 67.2325 49.688 69.3865 49.796 ;
          END
     END q[9]
     PIN ren
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 71.798 31.57 72.7035 31.626 ;
          END
     END ren
     PIN shutoff
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 77.244 31.57 78.1655 31.626 ;
          END
     END shutoff
     PIN sleep
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 79.4035 33.938 80.3265 33.994 ;
          END
     END sleep
     PIN wa[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 74.36 33.938 75.3245 33.994 ;
          END
     END wa[0]
     PIN wa[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 73.1475 33.938 74.178 33.994 ;
          END
     END wa[1]
     PIN wen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 73.262 31.57 74.15 31.626 ;
          END
     END wen
     PIN wpulse[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 75.887 30.004 77.144 30.08 ;
          END
     END wpulse[0]
     PIN wpulse[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 71.4065 29.28 72.45 29.356 ;
          END
     END wpulse[1]
     PIN wpulseen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 72.2125 30.004 73.099 30.08 ;
          END
     END wpulseen
     PIN clk
     DIRECTION input ;
          USE CLOCK ;
          PORT
               LAYER m4 ;
               RECT 69.8725 32.406 70.9045 32.462 ;
          END
     END clk
     PIN vddp
     SHAPE ABUTMENT ;
     DIRECTION input ;
          USE POWER ;
          PORT
               LAYER m4 ;
               RECT 0.48 0.958 63.049 1.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 1.846 57.036 1.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 10.678 63.049 10.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 11.566 57.036 11.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 12.298 63.049 12.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.186 57.036 13.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.918 63.049 13.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 14.806 57.036 14.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 15.538 63.049 15.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 16.426 57.036 16.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 17.158 63.049 17.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.046 57.036 18.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.778 63.049 18.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 19.666 57.036 19.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 2.578 63.049 2.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 20.398 63.049 20.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 21.286 57.036 21.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 22.018 63.049 22.094 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 22.906 57.036 22.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 23.638 63.049 23.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 24.526 57.036 24.602 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 25.258 63.049 25.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 26.146 57.036 26.222 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 3.466 57.036 3.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 39.478 63.049 39.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 4.198 63.049 4.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 40.366 57.036 40.442 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 41.098 63.049 41.174 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 41.986 57.036 42.062 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 42.718 63.049 42.794 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 43.606 57.036 43.682 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 44.338 63.049 44.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 45.226 57.036 45.302 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 45.958 63.049 46.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 46.846 57.036 46.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 47.578 63.049 47.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 48.466 57.036 48.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 49.198 63.049 49.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.086 57.036 5.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.818 63.049 5.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 50.086 57.036 50.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 50.818 63.049 50.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 51.706 57.036 51.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 52.438 63.049 52.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 53.326 57.036 53.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 54.058 63.049 54.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 54.946 57.036 55.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 55.678 63.049 55.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 56.566 57.036 56.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 57.298 63.049 57.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 58.186 57.036 58.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 58.918 63.049 58.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 59.806 57.036 59.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 6.706 57.036 6.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 60.538 63.049 60.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 61.426 57.036 61.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 62.158 63.049 62.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 63.046 57.036 63.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 63.778 63.049 63.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 64.666 57.036 64.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 7.438 63.049 7.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 8.326 57.036 8.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 9.058 63.049 9.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 9.946 57.036 10.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 28.028 57.208 28.104 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 28.588 137.884 28.664 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 28.984 137.884 29.06 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 29.28 57.208 29.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 30.004 57.208 30.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 31.072 56.56 31.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 31.57 57.208 31.626 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 32.406 57.208 32.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 33.324 56.56 33.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 34.336 137.884 34.412 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 35.06 137.884 35.136 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 35.356 137.884 35.432 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 35.752 137.884 35.828 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 36.312 137.884 36.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 38.256 137.884 38.364 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 26.644 81.252 26.72 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 26.776 81.252 26.852 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 27.04 60.613 27.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 27.896 81.252 27.972 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 28.456 61.0005 28.532 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 37.696 81.252 37.772 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 38.716 81.252 38.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.248 38.98 81.252 39.056 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.2565 33.938 61.2505 33.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.2565 34.204 60.8165 34.28 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.2565 34.632 60.5665 34.708 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.2565 35.62 60.5665 35.696 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.2565 35.884 60.5665 35.96 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.2565 37.004 60.5665 37.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.2565 37.3 60.5665 37.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.299 32.406 61.7495 32.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.302 31.57 62.0135 31.626 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.317 30.004 72.1325 30.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.38 29.28 61.212 29.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 1.08 75.3295 1.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 10.8 75.3295 10.876 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 12.42 75.3295 12.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 14.04 75.3295 14.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 15.66 75.3295 15.736 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 17.28 75.3295 17.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 18.9 75.3295 18.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 2.7 75.3295 2.776 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 20.52 75.3295 20.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 22.14 75.3295 22.216 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 23.76 75.3295 23.836 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 25.38 75.3295 25.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 39.6 75.3295 39.676 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 4.32 75.3295 4.396 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 41.22 75.3295 41.296 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 42.84 75.3295 42.916 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 44.46 75.3295 44.536 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 46.08 75.3295 46.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 47.7 75.3295 47.776 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 49.32 75.3295 49.396 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 5.94 75.3295 6.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 50.94 75.3295 51.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 52.56 75.3295 52.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 54.18 75.3295 54.256 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 55.8 75.3295 55.876 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 57.42 75.3295 57.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 59.04 75.3295 59.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 60.66 75.3295 60.736 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 62.28 75.3295 62.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 63.9 75.3295 63.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 7.56 75.3295 7.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 62.973 9.18 75.3295 9.256 ;
          END
          PORT
               LAYER m4 ;
               RECT 73.686 34.632 81.2055 34.688 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 0.958 138.02 1.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 10.678 138.02 10.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 12.298 138.02 12.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 13.918 138.02 13.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 15.538 138.02 15.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 17.158 138.02 17.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 18.778 138.02 18.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 2.578 138.02 2.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 20.398 138.02 20.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 22.018 138.02 22.094 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 23.638 138.02 23.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 25.258 138.02 25.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 39.478 138.02 39.554 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 4.198 138.02 4.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 41.098 138.02 41.174 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 42.718 138.02 42.794 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 44.338 138.02 44.414 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 45.958 138.02 46.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 47.578 138.02 47.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 49.198 138.02 49.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 5.818 138.02 5.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 50.818 138.02 50.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 52.438 138.02 52.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 54.058 138.02 54.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 55.678 138.02 55.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 57.298 138.02 57.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 58.918 138.02 58.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 60.538 138.02 60.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 62.158 138.02 62.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 63.778 138.02 63.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 7.438 138.02 7.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.2535 9.058 138.02 9.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 75.631 28.292 79.74 28.4 ;
          END
          PORT
               LAYER m4 ;
               RECT 76.4795 35.884 81.252 35.96 ;
          END
          PORT
               LAYER m4 ;
               RECT 76.6365 35.62 81.252 35.696 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.0775 37.004 81.252 37.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.3345 30.004 81.1125 30.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 77.859 29.28 81.252 29.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 78.0175 34.928 81.2525 35.004 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.292 28.028 137.884 28.104 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.292 30.004 137.884 30.08 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.292 31.57 137.884 31.626 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.292 32.406 137.884 32.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.332 29.28 137.884 29.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 1.846 138.02 1.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 11.566 138.02 11.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 13.186 138.02 13.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 14.806 138.02 14.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 16.426 138.02 16.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 18.046 138.02 18.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 19.666 138.02 19.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 21.286 138.02 21.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 22.906 138.02 22.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 24.526 138.02 24.602 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 26.146 138.02 26.222 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 3.466 138.02 3.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 40.366 138.02 40.442 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 41.986 138.02 42.062 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 43.606 138.02 43.682 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 45.226 138.02 45.302 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 46.846 138.02 46.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 48.466 138.02 48.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 5.086 138.02 5.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 50.086 138.02 50.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 51.706 138.02 51.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 53.326 138.02 53.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 54.946 138.02 55.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 56.566 138.02 56.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 58.186 138.02 58.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 59.806 138.02 59.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 6.706 138.02 6.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 61.426 138.02 61.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 63.046 138.02 63.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 64.666 138.02 64.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 8.326 138.02 8.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.397 9.946 138.02 10.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.94 31.072 137.884 31.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 81.94 33.324 137.884 33.368 ;
          END
     END vddp
     PIN vss
     SHAPE ABUTMENT ;
     DIRECTION inout ;
          USE GROUND ;
          PORT
               LAYER m4 ;
               RECT 0.48 0.592 138.02 0.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 10.312 138.02 10.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 11.932 138.02 12.008 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.552 138.02 13.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 15.172 138.02 15.248 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 16.792 138.02 16.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.412 138.02 18.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 2.212 138.02 2.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 20.032 138.02 20.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 21.652 138.02 21.728 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 23.272 138.02 23.348 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 24.892 138.02 24.968 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 26.512 138.02 26.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 3.832 138.02 3.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 39.112 138.02 39.188 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 40.732 138.02 40.808 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 42.352 138.02 42.428 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 43.972 138.02 44.048 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 45.592 138.02 45.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 47.212 138.02 47.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 48.832 138.02 48.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.452 138.02 5.528 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 50.452 138.02 50.528 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 52.072 138.02 52.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 53.692 138.02 53.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 55.312 138.02 55.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 56.932 138.02 57.008 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 58.552 138.02 58.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 60.172 138.02 60.248 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 61.792 138.02 61.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 63.412 138.02 63.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 65.032 138.02 65.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 7.072 138.02 7.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 8.692 138.02 8.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 27.172 81.94 27.28 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 27.468 81.94 27.576 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 29.544 81.94 29.652 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 30.566 57.208 30.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 30.982 81.94 31.026 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 32.08 81.94 32.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 33.414 81.94 33.458 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 33.83 57.208 33.874 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 34.764 81.94 34.872 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 36.84 81.94 36.948 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 37.136 81.94 37.244 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 37.96 81.94 38.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 38.552 81.94 38.66 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.3355 30.554 81.1275 30.61 ;
          END
          PORT
               LAYER m4 ;
               RECT 57.3665 33.836 81.2115 33.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 1.602 81.2155 1.678 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 11.322 81.2155 11.398 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 12.942 81.2155 13.018 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 14.562 81.2155 14.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 16.182 81.2155 16.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 17.802 81.2155 17.878 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 19.422 81.2155 19.498 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 21.042 81.2155 21.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 22.662 81.2155 22.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 24.282 81.2155 24.358 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 25.902 81.2155 25.978 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 3.222 81.2155 3.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 4.842 81.2155 4.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 40.122 81.2155 40.198 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 41.742 81.2155 41.818 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 43.362 81.2155 43.438 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 44.982 81.2155 45.058 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 46.602 81.2155 46.678 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 48.222 81.2155 48.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 49.842 81.2155 49.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 51.462 81.2155 51.538 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 53.082 81.2155 53.158 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 54.702 81.2155 54.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 56.322 81.2155 56.398 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 57.942 81.2155 58.018 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 59.562 81.2155 59.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 6.462 81.2155 6.538 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 61.182 81.2155 61.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 62.802 81.2155 62.878 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 64.422 81.2155 64.498 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 8.082 81.2155 8.158 ;
          END
          PORT
               LAYER m4 ;
               RECT 60.4615 9.702 81.2155 9.778 ;
          END
     END vss
     OBS
          LAYER m1 SPACING 0 ;
               RECT 0.248 0.198 138.252 65.502 ;
          LAYER m2 SPACING 0 ;
               RECT 0.32 0.268 138.18 65.432 ;
          LAYER m3 SPACING 0 ;
               RECT 0.342 0.24 138.158 65.46 ;
          LAYER m4 SPACING 0 ;
               RECT 0.32 0.31 138.18 65.34 ;
     END
END ip224uhdlp1p11rf_2048x32m4b2c1s0_t0r0p1d0a1m1h
END LIBRARY
