#############################################################################################
## Intel Confidential                                                                      ##
#############################################################################################
## Copyright 2022 Intel Corporation. The information contained herein is the proprietary   ##
## and confidential information of Intel or its licensors, and is supplied subject to, and ##
## may be used only in accordance with, previously executed agreements with Intel.         ##
## EXCEPT AS MAY OTHERWISE BE AGREED IN WRITING: (1) ALL MATERIALS FURNISHED BY INTEL      ##
## HEREUNDER ARE PROVIDED "AS IS" WITHOUT WARRANTY OF ANY KIND; (2) INTEL SPECIFICALLY     ##
## DISCLAIMS ANY WARRANTY OF NONINFRINGEMENT, FITNESS FOR A PARTICULAR PURPOSE OR          ##
## MERCHANTABILITY; AND (3) INTEL WILL NOT BE LIABLE FOR ANY COSTS OF PROCUREMENT OF       ##
## SUBSTITUTES, LOSS OF PROFITS, INTERRUPTION OF BUSINESS, OR FOR ANY OTHER SPECIAL,       ##
## CONSEQUENTIAL OR INCIDENTAL DAMAGES, HOWEVER CAUSED, WHETHER FOR BREACH OF WARRANTY,    ##
## CONTRACT, TORT, NEGLIGENCE, STRICT LIABILITY OR OTHERWISE.                              ##
#############################################################################################
#############################################################################################
##                                                                                         ##
##  Vendor:                Intel Corporation                                               ##
##  Product:               ip224uhdlp1p11rf                                                ##
##  Version:               r1.0.1                                                          ##
##  Technology:            p1222.4                                                         ##
##  Celltype:              MemoryIP                                                        ##
##  IP Owner:              Intel CMO                                                       ##
##  Creation Time:         Wed Sep 14 2022 15:16:16                                        ##
##  Memory Name:           ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p1d0a1m1h                  ##
##  Memory Name Generated: ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p1d0a1m1h                  ##
##                                                                                         ##
#############################################################################################

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
SITE ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p1d0a1m1h
  SIZE 83.204 by 117.54 ;
  SYMMETRY X Y ;
  CLASS CORE ;
END ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p1d0a1m1h


MACRO ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p1d0a1m1h
     FOREIGN ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p1d0a1m1h 0.00 0.00 ;
     ORIGIN 0.00 0.00 ;
     SIZE 83.204 by 117.54 ;
     SYMMETRY X Y ;
     CLASS BLOCK ;
     SITE ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p1d0a1m1h ;
     PIN adr[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 48.1595 62.924 49.3495 63 ;
          END
     END adr[0]
     PIN adr[10]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 35.707 62.924 36.837 63 ;
          END
     END adr[10]
     PIN adr[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 47.7645 61.804 48.7515 61.88 ;
          END
     END adr[1]
     PIN adr[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 34.4455 57.49 35.597 57.546 ;
          END
     END adr[2]
     PIN adr[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 47.59 60.848 48.764 60.924 ;
          END
     END adr[3]
     PIN adr[4]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 48.844 60.848 50.006 60.924 ;
          END
     END adr[4]
     PIN adr[5]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 33.045 52.96 34.002 53.036 ;
          END
     END adr[5]
     PIN adr[6]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 34.3265 58.326 35.266 58.382 ;
          END
     END adr[6]
     PIN adr[7]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 33.008 54.226 34.389 54.302 ;
          END
     END adr[7]
     PIN adr[8]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 33.4325 54.376 34.741 54.452 ;
          END
     END adr[8]
     PIN adr[9]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 35.695 61.804 36.6195 61.88 ;
          END
     END adr[9]
     PIN bc1
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 47.8445 61.54 48.9085 61.616 ;
          END
     END bc1
     PIN bc2
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 48.764 59.858 49.9035 59.914 ;
          END
     END bc2
     PIN clkbyp
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 44.767 58.326 45.6195 58.382 ;
          END
     END clkbyp
     PIN deepslp
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 49.268 58.326 50.262 58.382 ;
          END
     END deepslp
     PIN din[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 114.488 39.618 114.596 ;
          END
     END din[0]
     PIN din[10]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 82.088 39.618 82.196 ;
          END
     END din[10]
     PIN din[11]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 78.848 39.618 78.956 ;
          END
     END din[11]
     PIN din[12]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 75.608 39.618 75.716 ;
          END
     END din[12]
     PIN din[13]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 72.368 39.618 72.476 ;
          END
     END din[13]
     PIN din[14]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 69.128 39.618 69.236 ;
          END
     END din[14]
     PIN din[15]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 65.888 39.618 65.996 ;
          END
     END din[15]
     PIN din[16]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 50.048 39.618 50.156 ;
          END
     END din[16]
     PIN din[17]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 46.808 39.618 46.916 ;
          END
     END din[17]
     PIN din[18]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 43.568 39.618 43.676 ;
          END
     END din[18]
     PIN din[19]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 40.328 39.618 40.436 ;
          END
     END din[19]
     PIN din[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 111.248 39.618 111.356 ;
          END
     END din[1]
     PIN din[20]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 37.088 39.618 37.196 ;
          END
     END din[20]
     PIN din[21]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 33.848 39.618 33.956 ;
          END
     END din[21]
     PIN din[22]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 30.608 39.618 30.716 ;
          END
     END din[22]
     PIN din[23]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 27.368 39.618 27.476 ;
          END
     END din[23]
     PIN din[24]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 24.128 39.618 24.236 ;
          END
     END din[24]
     PIN din[25]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 20.888 39.618 20.996 ;
          END
     END din[25]
     PIN din[26]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 17.648 39.618 17.756 ;
          END
     END din[26]
     PIN din[27]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 14.408 39.618 14.516 ;
          END
     END din[27]
     PIN din[28]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 11.168 39.618 11.276 ;
          END
     END din[28]
     PIN din[29]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 7.928 39.618 8.036 ;
          END
     END din[29]
     PIN din[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 108.008 39.618 108.116 ;
          END
     END din[2]
     PIN din[30]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 4.688 39.618 4.796 ;
          END
     END din[30]
     PIN din[31]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 1.448 39.618 1.556 ;
          END
     END din[31]
     PIN din[3]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 104.768 39.618 104.876 ;
          END
     END din[3]
     PIN din[4]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 101.528 39.618 101.636 ;
          END
     END din[4]
     PIN din[5]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 98.288 39.618 98.396 ;
          END
     END din[5]
     PIN din[6]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 95.048 39.618 95.156 ;
          END
     END din[6]
     PIN din[7]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 91.808 39.618 91.916 ;
          END
     END din[7]
     PIN din[8]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 88.568 39.618 88.676 ;
          END
     END din[8]
     PIN din[9]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 36.766 85.328 39.618 85.436 ;
          END
     END din[9]
     PIN fwen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 48.4195 57.49 49.374 57.546 ;
          END
     END fwen
     PIN mc[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 35.244 60.124 36.283 60.2 ;
          END
     END mc[0]
     PIN mc[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 33.024 61.54 34.252 61.616 ;
          END
     END mc[1]
     PIN mc[2]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 34.383 61.54 35.525 61.616 ;
          END
     END mc[2]
     PIN mcen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 34.4805 61.804 35.417 61.88 ;
          END
     END mcen
     PIN mpr
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 47.125 57.49 48.061 57.546 ;
          END
     END mpr
     PIN q[0]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 114.488 41.423 114.596 ;
          END
     END q[0]
     PIN q[10]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 82.088 41.423 82.196 ;
          END
     END q[10]
     PIN q[11]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 78.848 41.423 78.956 ;
          END
     END q[11]
     PIN q[12]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 75.608 41.423 75.716 ;
          END
     END q[12]
     PIN q[13]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 72.368 41.423 72.476 ;
          END
     END q[13]
     PIN q[14]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 69.128 41.423 69.236 ;
          END
     END q[14]
     PIN q[15]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 65.888 41.423 65.996 ;
          END
     END q[15]
     PIN q[16]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 50.048 41.423 50.156 ;
          END
     END q[16]
     PIN q[17]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 46.808 41.423 46.916 ;
          END
     END q[17]
     PIN q[18]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 43.568 41.423 43.676 ;
          END
     END q[18]
     PIN q[19]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 40.328 41.423 40.436 ;
          END
     END q[19]
     PIN q[1]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 111.248 41.423 111.356 ;
          END
     END q[1]
     PIN q[20]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 37.088 41.423 37.196 ;
          END
     END q[20]
     PIN q[21]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 33.848 41.423 33.956 ;
          END
     END q[21]
     PIN q[22]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 30.608 41.423 30.716 ;
          END
     END q[22]
     PIN q[23]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 27.368 41.423 27.476 ;
          END
     END q[23]
     PIN q[24]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 24.128 41.423 24.236 ;
          END
     END q[24]
     PIN q[25]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 20.888 41.423 20.996 ;
          END
     END q[25]
     PIN q[26]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 17.648 41.423 17.756 ;
          END
     END q[26]
     PIN q[27]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 14.408 41.423 14.516 ;
          END
     END q[27]
     PIN q[28]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 11.168 41.423 11.276 ;
          END
     END q[28]
     PIN q[29]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 7.928 41.423 8.036 ;
          END
     END q[29]
     PIN q[2]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 108.008 41.423 108.116 ;
          END
     END q[2]
     PIN q[30]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 4.688 41.423 4.796 ;
          END
     END q[30]
     PIN q[31]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 1.448 41.423 1.556 ;
          END
     END q[31]
     PIN q[3]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 104.768 41.423 104.876 ;
          END
     END q[3]
     PIN q[4]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 101.528 41.423 101.636 ;
          END
     END q[4]
     PIN q[5]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 98.288 41.423 98.396 ;
          END
     END q[5]
     PIN q[6]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 95.048 41.423 95.156 ;
          END
     END q[6]
     PIN q[7]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 91.808 41.423 91.916 ;
          END
     END q[7]
     PIN q[8]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 88.568 41.423 88.676 ;
          END
     END q[8]
     PIN q[9]
     DIRECTION output ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 39.698 85.328 41.423 85.436 ;
          END
     END q[9]
     PIN ren
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 44.15 57.49 45.0555 57.546 ;
          END
     END ren
     PIN shutoff
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 49.596 57.49 50.5175 57.546 ;
          END
     END shutoff
     PIN sleep
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 51.7555 59.858 52.6785 59.914 ;
          END
     END sleep
     PIN wa[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 46.712 59.858 47.6765 59.914 ;
          END
     END wa[0]
     PIN wa[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 45.4995 59.858 46.53 59.914 ;
          END
     END wa[1]
     PIN wen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 45.614 57.49 46.502 57.546 ;
          END
     END wen
     PIN wpulse[0]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 48.239 55.924 49.496 56 ;
          END
     END wpulse[0]
     PIN wpulse[1]
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 43.7585 55.2 44.802 55.276 ;
          END
     END wpulse[1]
     PIN wpulseen
     DIRECTION input ;
          USE SIGNAL ;
          PORT
               LAYER m4 ;
               RECT 44.5645 55.924 45.451 56 ;
          END
     END wpulseen
     PIN clk
     DIRECTION input ;
          USE CLOCK ;
          PORT
               LAYER m4 ;
               RECT 42.2245 58.326 43.2565 58.382 ;
          END
     END clk
     PIN vddp
     SHAPE ABUTMENT ;
     DIRECTION input ;
          USE POWER ;
          PORT
               LAYER m4 ;
               RECT 0.48 0.958 35.401 1.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 1.846 29.388 1.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 10.678 35.401 10.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 100.306 29.388 100.382 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 101.038 35.401 101.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 101.926 29.388 102.002 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 102.658 35.487 102.734 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 103.546 29.388 103.622 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 104.278 35.401 104.354 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 105.166 29.388 105.242 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 105.898 35.487 105.974 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 106.786 29.388 106.862 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 107.518 35.401 107.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 108.406 29.388 108.482 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 109.138 35.487 109.214 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 11.566 29.388 11.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 110.026 29.388 110.102 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 110.758 35.401 110.834 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 111.646 29.388 111.722 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 112.378 35.487 112.454 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 113.266 29.388 113.342 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 113.998 35.401 114.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 114.886 29.388 114.962 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 115.618 35.487 115.694 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 116.506 29.388 116.582 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 12.298 35.487 12.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.186 29.388 13.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.918 35.401 13.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 14.806 29.388 14.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 15.538 35.487 15.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 16.426 29.388 16.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 17.158 35.401 17.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.046 29.388 18.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.778 35.487 18.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 19.666 29.388 19.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 2.578 35.487 2.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 20.398 35.401 20.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 21.286 29.388 21.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 22.018 35.487 22.094 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 22.906 29.388 22.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 23.638 35.401 23.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 24.526 29.388 24.602 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 25.258 35.487 25.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 26.146 29.388 26.222 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 26.878 35.401 26.954 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 27.766 29.388 27.842 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 28.498 35.487 28.574 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 29.386 29.388 29.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 3.466 29.388 3.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 30.118 35.401 30.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 31.006 29.388 31.082 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 31.738 35.487 31.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 32.626 29.388 32.702 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 33.358 35.401 33.434 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 34.246 29.388 34.322 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 34.978 35.487 35.054 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 35.866 29.388 35.942 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 36.598 35.401 36.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 37.486 29.388 37.562 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 38.218 35.487 38.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 39.106 29.388 39.182 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 39.838 35.401 39.914 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 4.198 35.401 4.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 40.726 29.388 40.802 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 41.458 35.487 41.534 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 42.346 29.388 42.422 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 43.078 35.401 43.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 43.966 29.388 44.042 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 44.698 35.487 44.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 45.586 29.388 45.662 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 46.318 35.401 46.394 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 47.206 29.388 47.282 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 47.938 35.487 48.014 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 48.826 29.388 48.902 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 49.558 35.401 49.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.086 29.388 5.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.818 35.487 5.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 50.446 29.388 50.522 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 51.178 35.487 51.254 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 52.066 29.388 52.142 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 6.706 29.388 6.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 65.398 35.401 65.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 66.286 29.388 66.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 67.018 35.487 67.094 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 67.906 29.388 67.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 68.638 35.401 68.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 69.526 29.388 69.602 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 7.438 35.401 7.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 70.258 35.487 70.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 71.146 29.388 71.222 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 71.878 35.401 71.954 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 72.766 29.388 72.842 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 73.498 35.487 73.574 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 74.386 29.388 74.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 75.118 35.401 75.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 76.006 29.388 76.082 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 76.738 35.487 76.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 77.626 29.388 77.702 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 78.358 35.401 78.434 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 79.246 29.388 79.322 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 79.978 35.487 80.054 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 8.326 29.388 8.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 80.866 29.388 80.942 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 81.598 35.401 81.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 82.486 29.388 82.562 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 83.218 35.487 83.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 84.106 29.388 84.182 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 84.838 35.401 84.914 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 85.726 29.388 85.802 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 86.458 35.487 86.534 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 87.346 29.388 87.422 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 88.078 35.401 88.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 88.966 29.388 89.042 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 89.698 35.487 89.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 9.058 35.487 9.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 9.946 29.388 10.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 90.586 29.388 90.662 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 91.318 35.401 91.394 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 92.206 29.388 92.282 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 92.938 35.487 93.014 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 93.826 29.388 93.902 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 94.558 35.401 94.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 95.446 29.388 95.522 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 96.178 35.487 96.254 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 97.066 29.388 97.142 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 97.798 35.401 97.874 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 98.686 29.388 98.762 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 99.418 35.487 99.494 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 53.948 29.56 54.024 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 54.508 82.588 54.584 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 54.904 82.588 54.98 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 55.2 29.56 55.276 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 55.924 29.56 56 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 56.992 28.912 57.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 57.49 29.56 57.546 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 58.326 29.56 58.382 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 59.244 28.912 59.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 60.256 82.588 60.332 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 60.98 82.588 61.056 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 61.276 82.588 61.352 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 61.672 82.588 61.748 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 62.232 82.588 62.308 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 64.176 82.588 64.284 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6 52.564 53.604 52.64 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6 52.696 53.604 52.772 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6 52.96 32.965 53.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6 53.816 53.604 53.892 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6 54.376 33.3525 54.452 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6 63.616 53.604 63.692 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6 64.636 53.604 64.712 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6 64.9 53.604 64.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6085 59.858 33.6025 59.914 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6085 60.124 33.1685 60.2 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6085 60.552 32.9185 60.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6085 61.54 32.9185 61.616 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6085 61.804 32.9185 61.88 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6085 62.924 32.9185 63 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6085 63.22 32.9185 63.296 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.651 58.326 34.1015 58.382 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.654 57.49 34.3655 57.546 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.669 55.924 44.4845 56 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.732 55.2 33.564 55.276 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 1.08 47.814 1.156 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 10.8 47.814 10.876 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 101.16 47.814 101.236 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 104.4 47.814 104.476 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 107.64 47.814 107.716 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 110.88 47.814 110.956 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 114.12 47.814 114.196 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 14.04 47.814 14.116 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 17.28 47.814 17.356 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 20.52 47.814 20.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 23.76 47.814 23.836 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 27 47.814 27.076 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 30.24 47.814 30.316 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 33.48 47.814 33.556 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 36.72 47.814 36.796 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 39.96 47.814 40.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 4.32 47.814 4.396 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 43.2 47.814 43.276 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 46.44 47.814 46.516 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 49.68 47.814 49.756 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 65.52 47.814 65.596 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 68.76 47.814 68.836 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 7.56 47.814 7.636 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 72 47.814 72.076 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 75.24 47.814 75.316 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 78.48 47.814 78.556 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 81.72 47.814 81.796 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 84.96 47.814 85.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 88.2 47.814 88.276 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 91.44 47.814 91.516 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 94.68 47.814 94.756 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.325 97.92 47.814 97.996 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 102.78 47.6575 102.856 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 106.02 47.6575 106.096 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 109.26 47.6575 109.336 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 112.5 47.6575 112.576 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 115.74 47.6575 115.816 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 12.42 47.6575 12.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 15.66 47.6575 15.736 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 18.9 47.6575 18.976 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 2.7 47.6575 2.776 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 22.14 47.6575 22.216 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 25.38 47.6575 25.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 28.62 47.6575 28.696 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 31.86 47.6575 31.936 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 35.1 47.6575 35.176 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 38.34 47.6575 38.416 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 41.58 47.6575 41.656 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 44.82 47.6575 44.896 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 48.06 47.6575 48.136 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 5.94 47.6575 6.016 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 51.3 47.6575 51.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 67.14 47.6575 67.216 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 70.38 47.6575 70.456 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 73.62 47.6575 73.696 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 76.86 47.6575 76.936 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 80.1 47.6575 80.176 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 83.34 47.6575 83.416 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 86.58 47.6575 86.656 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 89.82 47.6575 89.896 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 9.18 47.6575 9.256 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 93.06 47.6575 93.136 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 96.3 47.6575 96.376 ;
          END
          PORT
               LAYER m4 ;
               RECT 35.487 99.54 47.6575 99.616 ;
          END
          PORT
               LAYER m4 ;
               RECT 46.038 60.552 53.5575 60.608 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 102.658 82.724 102.734 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 105.898 82.724 105.974 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 109.138 82.724 109.214 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 112.378 82.724 112.454 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 115.618 82.724 115.694 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 12.298 82.724 12.374 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 15.538 82.724 15.614 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 18.778 82.724 18.854 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 2.578 82.724 2.654 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 22.018 82.724 22.094 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 25.258 82.724 25.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 28.498 82.724 28.574 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 31.738 82.724 31.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 34.978 82.724 35.054 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 38.218 82.724 38.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 41.458 82.724 41.534 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 44.698 82.724 44.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 47.938 82.724 48.014 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 5.818 82.724 5.894 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 51.178 82.724 51.254 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 67.018 82.724 67.094 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 70.258 82.724 70.334 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 73.498 82.724 73.574 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 76.738 82.724 76.814 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 79.978 82.724 80.054 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 83.218 82.724 83.294 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 86.458 82.724 86.534 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 89.698 82.724 89.774 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 9.058 82.724 9.134 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 92.938 82.724 93.014 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 96.178 82.724 96.254 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.5815 99.418 82.724 99.494 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 0.958 82.724 1.034 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 10.678 82.724 10.754 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 101.038 82.724 101.114 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 104.278 82.724 104.354 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 107.518 82.724 107.594 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 110.758 82.724 110.834 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 113.998 82.724 114.074 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 13.918 82.724 13.994 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 17.158 82.724 17.234 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 20.398 82.724 20.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 23.638 82.724 23.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 26.878 82.724 26.954 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 30.118 82.724 30.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 33.358 82.724 33.434 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 36.598 82.724 36.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 39.838 82.724 39.914 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 4.198 82.724 4.274 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 43.078 82.724 43.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 46.318 82.724 46.394 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 49.558 82.724 49.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 65.398 82.724 65.474 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 68.638 82.724 68.714 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 7.438 82.724 7.514 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 71.878 82.724 71.954 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 75.118 82.724 75.194 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 78.358 82.724 78.434 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 81.598 82.724 81.674 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 84.838 82.724 84.914 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 88.078 82.724 88.154 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 91.318 82.724 91.394 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 94.558 82.724 94.634 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.738 97.798 82.724 97.874 ;
          END
          PORT
               LAYER m4 ;
               RECT 47.983 54.212 52.092 54.32 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.8315 61.804 53.604 61.88 ;
          END
          PORT
               LAYER m4 ;
               RECT 48.9885 61.54 53.604 61.616 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.4295 62.924 53.604 63 ;
          END
          PORT
               LAYER m4 ;
               RECT 49.6865 55.924 53.4645 56 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.211 55.2 53.604 55.276 ;
          END
          PORT
               LAYER m4 ;
               RECT 50.3695 60.848 53.6045 60.924 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.644 53.948 82.588 54.024 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.644 55.924 82.588 56 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.644 57.49 82.588 57.546 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.644 58.326 82.588 58.382 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.684 55.2 82.588 55.276 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 1.846 82.724 1.922 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 100.306 82.724 100.382 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 101.926 82.724 102.002 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 103.546 82.724 103.622 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 105.166 82.724 105.242 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 106.786 82.724 106.862 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 108.406 82.724 108.482 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 11.566 82.724 11.642 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 110.026 82.724 110.102 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 111.646 82.724 111.722 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 113.266 82.724 113.342 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 114.886 82.724 114.962 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 116.506 82.724 116.582 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 13.186 82.724 13.262 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 14.806 82.724 14.882 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 16.426 82.724 16.502 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 18.046 82.724 18.122 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 19.666 82.724 19.742 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 21.286 82.724 21.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 22.906 82.724 22.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 24.526 82.724 24.602 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 26.146 82.724 26.222 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 27.766 82.724 27.842 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 29.386 82.724 29.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 3.466 82.724 3.542 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 31.006 82.724 31.082 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 32.626 82.724 32.702 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 34.246 82.724 34.322 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 35.866 82.724 35.942 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 37.486 82.724 37.562 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 39.106 82.724 39.182 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 40.726 82.724 40.802 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 42.346 82.724 42.422 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 43.966 82.724 44.042 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 45.586 82.724 45.662 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 47.206 82.724 47.282 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 48.826 82.724 48.902 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 5.086 82.724 5.162 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 50.446 82.724 50.522 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 52.066 82.724 52.142 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 6.706 82.724 6.782 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 66.286 82.724 66.362 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 67.906 82.724 67.982 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 69.526 82.724 69.602 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 71.146 82.724 71.222 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 72.766 82.724 72.842 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 74.386 82.724 74.462 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 76.006 82.724 76.082 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 77.626 82.724 77.702 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 79.246 82.724 79.322 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 8.326 82.724 8.402 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 80.866 82.724 80.942 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 82.486 82.724 82.562 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 84.106 82.724 84.182 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 85.726 82.724 85.802 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 87.346 82.724 87.422 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 88.966 82.724 89.042 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 9.946 82.724 10.022 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 90.586 82.724 90.662 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 92.206 82.724 92.282 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 93.826 82.724 93.902 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 95.446 82.724 95.522 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 97.066 82.724 97.142 ;
          END
          PORT
               LAYER m4 ;
               RECT 53.749 98.686 82.724 98.762 ;
          END
          PORT
               LAYER m4 ;
               RECT 54.292 56.992 82.588 57.036 ;
          END
          PORT
               LAYER m4 ;
               RECT 54.292 59.244 82.588 59.288 ;
          END
     END vddp
     PIN vss
     SHAPE ABUTMENT ;
     DIRECTION inout ;
          USE GROUND ;
          PORT
               LAYER m4 ;
               RECT 0.48 0.592 82.724 0.668 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 10.312 82.724 10.388 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 100.672 82.724 100.748 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 102.292 82.724 102.368 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 103.912 82.724 103.988 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 105.532 82.724 105.608 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 107.152 82.724 107.228 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 108.772 82.724 108.848 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 11.932 82.724 12.008 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 110.392 82.724 110.468 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 112.012 82.724 112.088 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 113.632 82.724 113.708 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 115.252 82.724 115.328 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 116.872 82.724 116.948 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 13.552 82.724 13.628 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 15.172 82.724 15.248 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 16.792 82.724 16.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 18.412 82.724 18.488 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 2.212 82.724 2.288 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 20.032 82.724 20.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 21.652 82.724 21.728 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 23.272 82.724 23.348 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 24.892 82.724 24.968 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 26.512 82.724 26.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 28.132 82.724 28.208 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 29.752 82.724 29.828 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 3.832 82.724 3.908 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 31.372 82.724 31.448 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 32.992 82.724 33.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 34.612 82.724 34.688 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 36.232 82.724 36.308 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 37.852 82.724 37.928 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 39.472 82.724 39.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 41.092 82.724 41.168 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 42.712 82.724 42.788 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 44.332 82.724 44.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 45.952 82.724 46.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 47.572 82.724 47.648 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 49.192 82.724 49.268 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 5.452 82.724 5.528 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 50.812 82.724 50.888 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 52.432 82.724 52.508 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 65.032 82.724 65.108 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 66.652 82.724 66.728 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 68.272 82.724 68.348 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 69.892 82.724 69.968 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 7.072 82.724 7.148 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 71.512 82.724 71.588 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 73.132 82.724 73.208 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 74.752 82.724 74.828 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 76.372 82.724 76.448 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 77.992 82.724 78.068 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 79.612 82.724 79.688 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 8.692 82.724 8.768 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 81.232 82.724 81.308 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 82.852 82.724 82.928 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 84.472 82.724 84.548 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 86.092 82.724 86.168 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 87.712 82.724 87.788 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 89.332 82.724 89.408 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 90.952 82.724 91.028 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 92.572 82.724 92.648 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 94.192 82.724 94.268 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 95.812 82.724 95.888 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 97.432 82.724 97.508 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.48 99.052 82.724 99.128 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 53.092 54.292 53.2 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 53.388 54.292 53.496 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 55.464 54.292 55.572 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 56.486 29.56 56.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 56.902 54.292 56.946 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 58 54.292 58.076 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 59.334 54.292 59.378 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 59.75 29.56 59.794 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 60.684 54.292 60.792 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 62.76 54.292 62.868 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 63.056 54.292 63.164 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 63.88 54.292 63.988 ;
          END
          PORT
               LAYER m4 ;
               RECT 0.616 64.472 54.292 64.58 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.6875 56.474 53.4795 56.53 ;
          END
          PORT
               LAYER m4 ;
               RECT 29.7185 59.756 53.5635 59.812 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 1.602 53.388 1.678 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 100.062 53.36 100.138 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 101.682 53.388 101.758 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 103.302 53.36 103.378 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 104.922 53.388 104.998 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 106.542 53.36 106.618 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 108.162 53.388 108.238 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 109.782 53.36 109.858 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 11.322 53.388 11.398 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 111.402 53.388 111.478 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 113.022 53.36 113.098 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 114.642 53.388 114.718 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 116.262 53.36 116.338 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 12.942 53.36 13.018 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 14.562 53.388 14.638 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 16.182 53.36 16.258 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 17.802 53.388 17.878 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 19.422 53.36 19.498 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 21.042 53.388 21.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 22.662 53.36 22.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 24.282 53.388 24.358 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 25.902 53.36 25.978 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 27.522 53.388 27.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 29.142 53.36 29.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 3.222 53.36 3.298 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 30.762 53.388 30.838 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 32.382 53.36 32.458 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 34.002 53.388 34.078 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 35.622 53.36 35.698 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 37.242 53.388 37.318 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 38.862 53.36 38.938 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 4.842 53.388 4.918 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 40.482 53.388 40.558 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 42.102 53.36 42.178 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 43.722 53.388 43.798 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 45.342 53.36 45.418 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 46.962 53.388 47.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 48.582 53.36 48.658 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 50.202 53.388 50.278 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 51.822 53.36 51.898 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 6.462 53.36 6.538 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 66.042 53.388 66.118 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 67.662 53.36 67.738 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 69.282 53.388 69.358 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 70.902 53.36 70.978 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 72.522 53.388 72.598 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 74.142 53.36 74.218 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 75.762 53.388 75.838 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 77.382 53.36 77.458 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 79.002 53.388 79.078 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 8.082 53.388 8.158 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 80.622 53.36 80.698 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 82.242 53.388 82.318 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 83.862 53.36 83.938 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 85.482 53.388 85.558 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 87.102 53.36 87.178 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 88.722 53.388 88.798 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 9.702 53.36 9.778 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 90.342 53.36 90.418 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 91.962 53.388 92.038 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 93.582 53.36 93.658 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 95.202 53.388 95.278 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 96.822 53.36 96.898 ;
          END
          PORT
               LAYER m4 ;
               RECT 32.8135 98.442 53.388 98.518 ;
          END
     END vss
     OBS
          LAYER m1 SPACING 0 ;
               RECT 0.248 0.198 82.956 117.342 ;
          LAYER m2 SPACING 0 ;
               RECT 0.32 0.268 82.884 117.272 ;
          LAYER m3 SPACING 0 ;
               RECT 0.342 0.24 82.862 117.3 ;
          LAYER m4 SPACING 0 ;
               RECT 0.32 0.31 82.884 117.18 ;
     END
END ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p1d0a1m1h
END LIBRARY
